module main;
initial
begin
$display("goodbye world");
$finish;
end
endmodule
